interface intf(input logic rst);
  
  logic [7:0] a;
  logic [7:0] b;
  logic [7:0] c;
  logic [7:0] sum;
  logic [1:0] carry;
  
endinterface: intf